library IEEE;
use IEEE.std_logic_1164.all;

--Figure out how to create a 2D array of components. 
entity Systolic is 
    port(load, clr, clk: in std_logic);
end Systolic;